library IEEE; 
use IEEE.std_logic_1164.all;

package int_array is 

type array_of_int_5 is array (0 to 4) of integer;

end int_array;
