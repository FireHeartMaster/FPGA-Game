library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity character_rom2 is
  
  port (
    addr : in  unsigned(8 downto 0);
    clk  : in  std_logic;
    dout : out unsigned(3 downto 0));
end character_rom2;

architecture rtl of character_rom2 is
  type rom_array is array (0 to 399) of unsigned(3 downto 0);

  constant ROM : rom_array := (
   "0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0100",
	"0010",
	"0001",
	"0001",
	"0010",
	"0100",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0010",
	"0100",
	"0111",
	"1001",
	"1011",
	"1011",
	"1001",
	"0111",
	"0100",
	"0010",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0011",
	"0101",
	"1010",
	"1110",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1110",
	"1010",
	"0101",
	"0011",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0010",
	"0110",
	"1101",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1101",
	"0110",
	"0010",
	"0000",
	"0000",
	"0000",
	"0011",
	"0101",
	"1101",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1110",
	"0110",
	"0011",
	"0000",
	"0000",
	"0010",
	"1011",
	"1111",
	"1110",
	"1101",
	"1110",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1110",
	"1101",
	"1110",
	"1111",
	"1011",
	"0010",
	"0000",
	"0011",
	"0100",
	"1110",
	"1001",
	"0101",
	"0010",
	"0110",
	"1100",
	"1111",
	"1111",
	"1111",
	"1111",
	"1100",
	"0111",
	"0011",
	"0100",
	"1000",
	"1110",
	"0100",
	"0011",
	"0001",
	"0101",
	"1100",
	"1000",
	"1001",
	"0010",
	"0011",
	"0111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1001",
	"1011",
	"0101",
	"0001",
	"0011",
	"1100",
	"0101",
	"0001",
	"0001",
	"0101",
	"1100",
	"0101",
	"0011",
	"0001",
	"0100",
	"1001",
	"1111",
	"1111",
	"1111",
	"1111",
	"1000",
	"0100",
	"0010",
	"0011",
	"0110",
	"1100",
	"0110",
	"0001",
	"0001",
	"0101",
	"1110",
	"1010",
	"0110",
	"0101",
	"1000",
	"1100",
	"1101",
	"1101",
	"1101",
	"1101",
	"1100",
	"1000",
	"0101",
	"0110",
	"1010",
	"1110",
	"0110",
	"0001",
	"0001",
	"0101",
	"1101",
	"1100",
	"1110",
	"1111",
	"1111",
	"0111",
	"0010",
	"0011",
	"0011",
	"0010",
	"0111",
	"1111",
	"1110",
	"1110",
	"1100",
	"1101",
	"0110",
	"0001",
	"0001",
	"0101",
	"1110",
	"1101",
	"1111",
	"1111",
	"1111",
	"1001",
	"0011",
	"0100",
	"0100",
	"0011",
	"1000",
	"1111",
	"1111",
	"1111",
	"1101",
	"1110",
	"0110",
	"0001",
	"0001",
	"0101",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1110",
	"1001",
	"0110",
	"0110",
	"1001",
	"1110",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"0110",
	"0001",
	"0001",
	"0101",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1101",
	"1101",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"0110",
	"0000",
	"0000",
	"0101",
	"1011",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1111",
	"1011",
	"0000",
	"0000",
	"1011",
	"1011",
	"1111",
	"1111",
	"1011",
	"1011",
	"1111",
	"1111",
	"1111",
	"1111",
	"1001",
	"1001",
	"1111",
	"1111",
	"1111",
	"1111",
	"1010",
	"1011",
	"0000",
	"0000",
	"0010",
	"0001",
	"1011",
	"1011",
	"0010",
	"0010",
	"1001",
	"1111",
	"1111",
	"1001",
	"0010",
	"0001",
	"1000",
	"1111",
	"1111",
	"1001",
	"0010",
	"0010",
	"0000",
	"0000",
	"0000",
	"0001",
	"1000",
	"1000",
	"0000",
	"0000",
	"0001",
	"1000",
	"1000",
	"0001",
	"0000",
	"0000",
	"0001",
	"1000",
	"1000",
	"0001",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0001",
	"0001",
	"0000",
	"0000",
	"0000",
	"0000",
	"0001",
	"0001",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000",
	"0000");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      dout <= ROM(TO_INTEGER(addr));
    end if;
  end process;

end rtl;
