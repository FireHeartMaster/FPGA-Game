library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity block_rom is
  
  port (
    addr : in  unsigned(8 downto 0);
    clk  : in  std_logic;
    dout : out unsigned(3 downto 0));
end block_rom;

architecture rtl of block_rom is
  type rom_array is array (0 to 399) of unsigned(3 downto 0);

  constant ROM : rom_array := (
   "0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0101",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0100",
	"0101",
	"0100",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0101",
	"0100",
	"0100",
	"0101",
	"0101");

begin

  process (clk)
  begin
    if rising_edge(clk) then
      dout <= ROM(TO_INTEGER(addr));
    end if;
  end process;

end rtl;
